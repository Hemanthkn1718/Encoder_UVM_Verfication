package en_pkg;

	import uvm_pkg::*;
	`include "uvm_macros.svh"

	`include "wr_cfg.sv"
	`include "rd_cfg.sv"
	`include "env_config.sv"

	`include "wr_xtn.sv"
	`include "wr_driver.sv"
	`include "wr_monitor.sv"
	`include "wr_sequencer.sv"
	`include "wr_seqs.sv"
	`include "wr_agent.sv"
	`include "wr_agent_top.sv"

	`include "rd_xtn.sv"
	`include "rd_driver.sv"
        `include "rd_monitor.sv"
        `include "rd_sequencer.sv"
        `include "rd_agent.sv"
        `include "rd_agent_top.sv"

 	`include "scoreboard.sv"
	`include "env.sv"
	`include "test.sv"
endpackage
